package test_pkg;
`include "msg_seq_item.sv"
`include "msg_seq.sv"
`include "msg_driver.sv"
`include "msg_monitor.sv"
`include "msg_agent.sv"
// `include "sim/uvm/hash_if.sv"
`include "hash_seq_item.sv"
`include "hash_seq.sv"
`include "hash_driver.sv"
`include "hash_monitor.sv"
`include "hash_agent.sv"
`include "sha_scoreboard.sv"
`include "sha_env.sv"
// `include "src/rtl/sha_algo_wrapper.sv"
// `include "sim/sha_uvm_tb_top.sv"
// `include "sim/single_value_test.sv"

endpackage // test_pkg
   
